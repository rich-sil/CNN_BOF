library IEEE, STD;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.FIXED_PKG.ALL;
use STD.TEXTIO.ALL;

entity conv_4 is
    Port ( clk : in STD_LOGIC;
           ready_in : in STD_LOGIC;
           in_4 : in STD_LOGIC_VECTOR (191 downto 0);
           start_out : out STD_LOGIC := '0';
           last_out : out STD_LOGIC := '0';
           pop_out : out STD_LOGIC := '0';
           conv4_out : out STD_LOGIC_VECTOR (399 downto 0) );
end conv_4; 

architecture Behavioral of conv_4 is

constant int : INTEGER := 1;
constant dec : INTEGER := -7;

constant int_2 : INTEGER := 3;
constant dec_2 : INTEGER := -12;

constant int_buff : INTEGER := 3;
constant dec_buff : INTEGER := -12;

constant up : INTEGER := 191;
constant down : INTEGER := 176;
constant bits : INTEGER := 16;

type w is array (0 to 1499) of sfixed (int downto dec);
signal weights : w :=     (
                            "000000000", "000000000", "111100110", "111110101", "111001100", "000000110", "111000010", "111110001", "000010101", "000001111", 
                            "110110111", "000011000", "111011000", "111110101", "000000001", "111010111", "111100100", "111110101", "111000010", "111111001", 
                            "111111001", "000010000", "000000011", "111101110", "110110100", "000010010", "000000111", "111010110", "111010010", "000111010", 
                            "110110011", "000001011", "111101111", "111111011", "000000101", "000010100", "111001101", "000010011", "000011011", "111100001", 
                            "000011101", "000001100", "110110100", "111110101", "000010011", "000011011", "000111010", "001000001", "111111100", "000101001", 
                            "000011110", "111111110", "000100000", "000101100", "110111010", "111110100", "111110111", "111110000", "001000110", "001010010", 
                            "111100010", "000011100", "110111100", "111100000", "111100011", "000000101", "111100011", "000001011", "111110111", "000010011", "000010000", "111001111", "000001101", "000001110", "110000011", "000000001", "000000101", "110110101", "000010011", "111111101", "111111110", "000010000", "111111011", "111001011", "000101011", "111101110", "111110010", "000101101", "111110100", "110011100", "000110100", "111101100", "000001101", "000001011", "111000001", "111010001", "000011110", "110111000", "001000001", "000010100", "111110110", "110110100", "000101110", "000100101", "111101110", "000000101", "110101111", "000111101", "000110001", "110110110", "001010100", "111100010", "111101010", "000001101", "000110110", "000100010", "000000001", "000001010", "111000000", "000110110", "110110010", "111100110", "110111000", "111110101", "111011011", "111010100", "111100111", "111111010", "000000011", "000000110", "111111101", "111100100", "111110011", "000000010", "000001101", "000010100", "000001001", "000000000", "000011010", "111110101", "000000110", "111101010", "000010101", "000001011", "000010101", "111111110", "111111101", "000000110", "000011001", "111101011", "110111001", "111011101", "000000100", "111101110", "000011010", "111111001", "111100110", "000001111", "000100000", "111111100", "111110011", "000101011", "111110111", "111111110", "000010101", "111110111", "000010100", "111110010", "000001010", "111110101", "000000000", "000110111", "000100001", "000100010", "001110100", "000010001", "000001010", "000010000", "111100110", "110100111", "111111100", "111110000", "111111000", "111111010", "000000101", "000000001", "111101110", "000010000", "111111011", "111110001", "000000100", "111110101", "111111110", "000000011", "111110001", "111111010", "000001010", "111101110", "000000111", "000001110", "000010000", "000000101", "111101111", "000000000", "111100100", "111101001", "111101111", "111101000", "000001101", "111110000", "111100111", "000001110", "000000111", "000000010", "111110101", "000000101", "111101001", "111110110", "111111000", "000001100", "000001110", "111101100", "111101110", "111101010", "111110110", "000001001", "000000010", "111110100", "000000110", "000000101", "000001001", "111101100", "111100110", "111100101", "000001101", "111111011", "111111000", "000000111", "111110000", "000000000", "111111111", "111101100", "000000110", "111111111", 
                            "111100110", "111111101", "111101001", "000000101", "000001110", "000010110", "000000001", "111111101", "111111100", "111110111", "111100100", "000000101", "111101111", "111101000", "111111000", "000010000", "000001101", "000000101", "000001010", "000010011", "111101001", "111111001", "000001001", "111110110", "000000100", "111101101", "111111111", "111110001", "000000000", "111111110", "111110001", "111111111", "111111111", "000000100", "000001101", "000000000", "111110100", "111111100", "111110111", "000010101", "000010010", "111101010", "111100111", "111101101", "000001101", "000001101", "111110011", "000001110", "111100111", "111111100", "000010010", "111111100", "000010110", "111101101", "000010011", "000000011", "111011010", "000011110", "000010100", "111101100", "111110001", "000001111", "000001110", "000010110", "000000100", "000000000", "000010111", "000100111", "111110111", "111111100", "111001101", "000111100", "000011110", "000010111", "001011110", "000000100", "111101010", "000000000", "111111010", "111011001", "000000000", "000001011", "010100100", "111000111", "111010101", "000101100", "110111000", "000010010", "111110001", "000001011", "111101111", "001011000", "111111011", "111101010", "111011100", "000010110", "000001101", "000100010", "000001101", "000100001", "000000001", "000000101", "111111000", "111010001", "111011111", "111100010", "000000000", "000011000", "000010100", "000000001", "000100101", "111111110", "111101111", "000000111", "111110000", "000010011", "111001010", "111111010", "110011001", "000011000", "001000000", "001010000", "000111001", "111111100", "000000100", "111111000", "111110010", "111100010", "000011010", "111111100", "010001110", "111100110", "111101100", "001000100", "111010111", "111101111", "111101110", "000001010", "111110100", "001111110", "000011111", "000010001", "111100111", "111100101", "000010001", "111101100", "111001001", "000000010", "111110000", "111111000", "000010100", "111101100", "111101000", "111111011", "111100000", "000101010", "111110011", "111110100", "111100000", "000000000", "000001011", "111101110", "111110101", "111000001", "111100101", "000000000", "001011001", "111111011", "000000011", "000000000", "111001100", "111111010", "000000101", "000000100", "000011011", "000001100", "111101111", "111110011", "000000101", "111111010", "000001011", "111111001", "000010000", "111110100", "000001111", "000001010", "111110000", "000010011", "111110100", "111101100", "000001011", "111110110", "111111100", "111111100", "000001101", "111101011", "111110000", "000001010", "111111101", "000001100", "111101000", "111110100", "111101101", "111111010", "000000110", "000000001", "000010001", "000000001", "000001010", "111111100", "111110011", "111110001", "000001001", "111111101", "111101010", "000000101", "111111100", "111101000", "000001111", "000001111", "111101110", "000001011", "000000000", "111110110", "111101001", "111110001", "111111110", "000001100", "111100111", "111110010", "111101100", "000001000", "000001010", "111110111", "111110011", "000000100", "000111101", "111010111", "001001101", "111111100", "111011101", "000011111", "111111110", "000001011", 
                            "000001101", "000010010", "111101111", "000100111", "111111100", "000000011", "000001011", "111011111", "111011101", "000011010", "111010111", "111011011", "111111011", "111111011", "111101111", "000110000", "111111011", "000010010", "000000001", "111010100", "000001001", "000000010", "110100011", "000000011", "111110001", "000001100", "000010111", "000000100", "111110010", "111111011", "110111010", "111110001", "111111010", "111101010", "110010100", "111111111", "111110000", "111110011", "000011000", "111110101", "111010110", "000011001", "110110011", "000100111", "000000101", "000100011", "000001000", "000100011", "000001101", "000010001", "000100110", "110011000", "110110111", "000011100", "111011110", "000100001", "000011101", "000001101", "111101101", "111111111", "111111100", "111111000", "000001010", "000011011", "111110010", "000001111", "111001101", "000101010", "000100110", "000001011", "000110111", "111101000", "111110100", "111111001", "111100001", "110011010", "000010101", "000001101", "000000100", "000001101", "111110100", "111011101", "000100000", "000010000", "111111011", "111111010", "111001100", "111111111", "111110110", "111100111", "111100100", "111000101", "111000101", "111100111", "111010101", "000001000", "111111110", "111110101", "000000000", "000100010", "110101011", "111111110", "000110011", "111001101", "111111101", "001001111", "111000111", "000000010", "000000110", "111101011", "000100111", "000101111", "000010100", "000011100", "001001000", "000001001", "000101100", "110101011", "000111011", "000001111", "111111100", "000010101", "000110011", "110111110", "000000001", "000000100", "000011110", "000011010", "000100011", "111001011", "000100111", "111110100", "000000100", "111111111", "111111010", "110001010", "111111011", "000001110", "000011011", "111011110", "111100100", "111110111", "000000111", "111110001", "111101010", "111110000", "111101100", "111010110", "000001010", "111101001", "111101100", "000010011", "111100111", "111101110", "000000001", "111100110", "111110111", "000010011", "111010110", "111011110", "000010110", "111011111", "111100011", "000001100", "111110000", "111001111", "000101111", "000001010", "000000011", "000000011", "111001110", "110110100", "000101111", "111110001", "000101110", "000000110", "111111010", "000000110", "000110100", "000001110", "111101100", "000000101", "111110010", "111101101", "000000010", "111101011", "000010000", "111110010", "111101111", "111111010", "000000101", "000100010", "111101100", "000001100", "111011100", "000000110", "111011101", "111111101", "000100000", "111100010", "000000000", "000010001", "111001000", "000000111", "111110110", "111110010", "000101000", "000100010", "000000100", "111111101", "000011001", "000010001", "000100110", "000001010", "000100111", "000000001", "111110101", "111111001", "000001001", "111110100", "000001000", "000001000", "000100001", "000100110", "000010111", "111111001", "000011001", "000010000", "000000100", "000000111", "111100010", "000001000", "111111110", "000001011", "111111100", "000010110", "111111001", "111010001", "111010000", "111100101", "111111100", "111110010", "000010100", "111101000", 
                            "111101111", "000011001", "110111010", "000000011", "111110101", "111001011", "111101100", "111111011", "111111110", "000010000", "000010001", "111010111", "111111010", "000010100", "111001110", "111100010", "000010001", "111101010", "111110110", "000000100", "000010010", "111110111", "000001000", "111111000", "111111000", "000001111", "111100100", "000000000", "000001011", "000111011", "111101001", "111110011", "111111000", "111110011", "111111001", "000010010", "111111101", "000011011", "000010010", "000001101", "000001001", "111110101", "000110000", "111100101", "000001101", "111101010", "000010110", "111101110", "111110110", "000011100", "111001111", "000010111", "000001110", "111101110", "111011100", "111111011", "111111010", "000000111", "000001110", "000000101", "111010100", "000000000", "000000100", "000010010", "111110110", "000010001", "111111110", "111110111", "000010101", "111111000", "000010011", "000010100", "111011111", "000001001", "000101001", "000000000", "000100000", "000001101", "111011101", "000001001", "111110011", "000000111", "000100101", "111110010", "111100010", "000011101", "111101001", "111101110", "000001101", "000001110", "111000011", "111100111", "111101111", "111110101", "000011111", "111110101", "111010011", "000000110", "111011100", "111100101", "000000111", "111111000", "111001110", "111101100", "111101010", "000000011", "000001100", "111110101", "000110011", "000000010", "001111111", "111100011", "111101010", "000101100", "111100100", "000001000", "111111000", "000010011", "111101110", "000101110", "111101111", "111111011", "110111111", "110111011", "111110011", "000010001", "111101010", "000011001", "111110110", "111111000", "000011101", "000111011", "111110010", "111111000", "111110101", "000111100", "000011110", "111101001", "000101111", "111111000", "000000010", "111111001", "000010100", "111010100", "000010101", "000000001", "000011110", "000011100", "000010100", "110110011", "111111100", "111010011", "000000110", "111110010", "111100110", "111101100", "111100000", "000011100", "111110110", "110110101", "111000001", "111111110", "110100011", "111101110", "000000101", "000010010", "000011011", "001001100", "110010110", "111110100", "111000110", "111011111", "111011110", "000101101", "111001101", "111110110", "000010010", "111101010", "000100100", "001101101", "000000011", "111101010", "000100000", "000010011", "000011110", "000011101", "000000010", "111111101", "111111011", "111111100", "000010011", "111110111", "000000010", "000010011", "000010111", "000011111", "000010100", "000010100", "000011110", "000010100", "000010001", "000000001", "000001100", "111011011", "000010111", "111100110", "000000101", "000100010", "000010100", "111101011", "000111110", "111111110", "111101110", "000000011", "111101001", "101111101", "000001010", "111011101", "000100101", "111011100", "111110100", "111100001", "000000010", "000000001", "000001000", "000010101", "111100000", "111010111", "111110001", "000000100", "111101111", "111101000", "000001101", "111111100", "111101011", "000000001", "111110010", "111111001", "111110100", "111101100", "000001010", "000000010", "000000000", "111111101", 
                            "000000110", "111100101", "000001111", "000010000", "111110110", "111111111", "111111111", "111111110", "111101110", "111100111", "000001010", "111110001", "111110100", "111110000", "000000011", "111110001", "111101101", "000000000", "111101001", "000001010", "000001100", "000000010", "000000011", "111101001", "000001001", "111111000", "000001000", "111110011", "000001100", "000000100", "111101101", "000001100", "000001010", "111110111", "111100101", "000001101", "111101010", "000000101", "000001011", "111111110", "111101100", "000001011", "111101011", "111101000", "111110000", "111111100", "110011000", "000001101", "000010011", "111000010", "111101011", "111101100", "000000010", "000010000", "000101001", "110010111", "111011011", "000011010", "110011001", "111111110", "000001011", "111011010", "111110001", "111111110", "000001110", "000000111", "111111001", "110110000", "000011001", "000000110", "110001010", "000010111", "000001111", "000000000", "111101000", "000000001", "000001101", "000000011", "000100001", "000001001", "000000010", "000011110", "111101110", "000101000", "000001111", "111110110", "000110000", "000000110", "111101111", "000010110", "111111101", "111001111", "000000100", "111111100", "111101100", "111111101", "000100001", "111000010", "000110110", "000010101", "000001111", "111111010", "111101111", "111011011", "000001010", "000000001", "000001101", "000001100", "000001000", "111110110", "111100111", "111111110", "111101010", "000010110", "000001001", "000000010", "111101111", "111101001", "000010011", "111100110", "111101010", "111111111", "111111001", "000000000", "111110001", "000010011", "111100110", "000001011", "000000000", "111110010", "111111111", "111111111", "000001110", "111101100", "111111110", "000000001", "000000010", "111110100", "111110111", "111110011", "000000100", "111111000", "111100011", "111110000", "000001110", "111110111", "111101001", "000010001", "000000010", "111110111", "000010000", "000001010", "111110101", "111101110", "000001100", "000001111", "111110001", "111110101", "000001001", "000001010", "111101010", "111101010", "111110100", "111101011", "000011010", "111101101", "111101001", "000011111", "000011111", "110101111", "000110101", "000000001", "111110010", "000010010", "111011000", "101000001", "000110001", "110000001", "000100100", "000100101", "000000101", "111000111", "000111111", "000000011", "111101011", "000001010", "101110001", "001101001", "000110011", "110001100", "001010011", "111010011", "110100100", "001000110", "000110110", "000101100", "000000000", "111110001", "111011000", "001101000", "111110000", "101111101", "001101011", "101010011", "111010111", "000110100", "000101010", "000101010", "000000101", "111111010", "111100100", "001001011", "111000101", "110111010", "000110100", "101011101", "111000100", "000111011", "110101100", "000101011", "000000000", "111101111", "111001100", "000011010", "000001101", "111110000", "000000100", "111101101", "111101001", "111101101", "111101101", "111111001", "000001110", "111101100", "111111000", "111111110", "111110011", "000010001", "111111000", "000000111", "000000000", "111111011", "111111000", "000001110", 
                            "000000010", "000001001", "111111000", "000000011", "000000001", "111110001", "000000001", "111110111", "000000010", "111111110", "000000010", "111111100", "111101100", "111111011", "111111100", "111111011", "000001011", "111111101", "111110101", "111101100", "000000000", "111111000", "000001110", "000000111", "000001111", "000001100", "000010010", "000001010", "000001010", "111111011", "111110001", "111110011", "111101000", "111110011", "000000000", "000001001", "111110111", "111111011", "111110010", "111101111", "111111101", "000001101", "000010010", "111110100", "000000001", "111110111", "111110101", "111110010", "111110000", "000001101", "000010100", "000010001", "000001001", "111100101", "111111010", "111101111", "111111000", "111101001", "000000000", "000000100", "000000110", "111101010", "111101011", "111111001", "111111011", "000000011", "111110010", "111111110", "000000101", "111110001", "000001000", "111111100", "000000110", "111111011", "000001010", "111111111", "111110010", "000000110", "111111010", "111111010", "111101110", "111100010", "000010110", "111110110", "000001101", "000001010", "111111100", "111111100", "111111001", "111110001", "000000001", "111111000", "000001010", "111101101", "000000011", "000010011", "111110011", "111111011", "111100110", "111110110", "000001001", "111100110", "000100110", "111101001", "111000101", "111100110", "000100001", "000000000", "111110100", "000001100", "111111101", "000110011", "000001010", "111110011", "000100000", "111100111", "111100101", "000100010", "111110001", "111110001", "000000001", "111111110", "000001000", "001000110", "000000111", "111111001", "000001111", "000110010", "000011011", "000100100", "000011101", "111111111", "111101110", "000010010", "000001000", "111100100", "000011011", "111011000", "000010011", "000010010", "111111011", "110111011", "000111000", "000000000", "000000000", "000010101", "111011100", "110100000", "000011111", "111010111", "111101110", "111111000", "111101100", "111011001", "000001101", "000100010", "000001001", "111110010", "111000010", "111011111", "111101001", "111100111", "111101101", "000001010", "111101011", "111110111", "111110000", "000000000", "000001100", "000001010", "111101001", "000010011", "111101010", "111101000", "111111011", "111110000", "111101110", "000010011", "000010011", "111101011", "111101111", "000010000", "111111010", "111101100", "111111011", "111110111", "111110000", "000001011", "000001110", "000000000", "000001110", "111111010", "000001110", "000000000", "000000100", "000001100", "111110110", "000010001", "000000101", "000001100", "000000011", "000000100", "000000000", "111111101", "111110001", "111111011", "111110001", "111110110", "111110100", "111101111", "000001100", "000000000", "000000000", "000001110", "111101100", "111110001", "111110001", "000010000", "111110011", "000000010", "111010000", "111111011", "000010100", "000011110", "000101000", "000001100", "000100000", "000011100", "111101011", "111110010", "000101011", "000011100", "111110101", "000000010", "001000001", "111111000", "000011100", "001010010", "000101000", "000110100", "111111110", "000010110", "111111001", "001000010", 
                            "000001000", "111110011", "000100110", "000011000", "000000000", "000111011", "000011010", "111110010", "111101111", "000000001", "111111001", "110100001", "000010010", "111010111", "000100110", "111111000", "111011111", "000010010", "000001010", "000011001", "111110010", "111111000", "110110110", "000000000", "000001010", "111010101", "000000111", "111110100", "111001100", "000001111", "111111111", "000000001", "111101111", "000001001", "111010110", "111001110" );
                            
type b is array (0 to 24) of sfixed (int downto dec);
signal bias : b :=        ( "111110001", "111101110", "111111101", "111111100", "111111101", "111001100", "111010110", "111111101", 
                            "000001100", "000001000", "000101111", "111110000", "000000110", "111110111", "111100101", "111111101", 
                            "111111011", "000001111", "111111010", "110101100", "111111011", "111111100", "000010110", "111111101", 
                            "000000111" );

type buff is array (0 to 24) of sfixed (int_buff downto dec_buff);
signal buff_1 : buff :=     ( others => X"0000" );

signal aux : UNSIGNED (2 downto 0) := "000";
signal cont : UNSIGNED (4 downto 0) := "00000";
signal k_cont : UNSIGNED (4 downto 0) := "00000";
signal temp : STD_LOGIC_VECTOR (up downto 0);
constant zero_out : STD_LOGIC_VECTOR := X"0000";

--constant int_out : INTEGER := 2;
--constant dec_out : INTEGER := -13;
--type p is array (0 to 11) of STD_LOGIC_VECTOR (8 downto 0);
--signal pesos : p :=     ( others => "000000000" );

--type m is array (0 to 11) of sfixed (int_2 downto dec_2);
--signal mults : m :=     ( others => X"0000");

--type res is array (0 to 24) of sfixed (15 downto -16);
--signal resultado : res :=   (others =>  X"00000000");
        
begin

    process(clk, ready_in, in_4)
    begin
    
        if rising_edge(clk) then
        
            if ( ready_in = '1' ) then
            
                if ( cont < 15 ) then
                    
                    if ( k_cont = 0 ) then
                    
                        pop_out <= '1';
                        start_out <= '0';
                        k_cont <= k_cont + 1;
                        
                        if ( aux = 4 ) then
                        
                            buff_1(to_integer(k_cont)) <= resize (  to_sfixed(in_4(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)) +
                                                                    to_sfixed(in_4(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1) +
                                                                    to_sfixed(in_4(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2) +
                                                                    to_sfixed(in_4(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3) + 
                                                                    to_sfixed(in_4(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4) +
                                                                    to_sfixed(in_4(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5) +
                                                                    to_sfixed(in_4(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6) +
                                                                    to_sfixed(in_4(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7) +
                                                                    to_sfixed(in_4(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8) +
                                                                    to_sfixed(in_4(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9) +
                                                                    to_sfixed(in_4(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10) +
                                                                    to_sfixed(in_4(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11) + 
                                                                    buff_1(to_integer(k_cont)) + bias(0), int_buff, dec_buff, fixed_saturate, fixed_truncate );                                                                    
                        else
                        
                            buff_1(to_integer(k_cont)) <= resize (  to_sfixed(in_4(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)) +
                                                                    to_sfixed(in_4(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1) +
                                                                    to_sfixed(in_4(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2) +
                                                                    to_sfixed(in_4(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3) + 
                                                                    to_sfixed(in_4(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4) +
                                                                    to_sfixed(in_4(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5) +
                                                                    to_sfixed(in_4(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6) +
                                                                    to_sfixed(in_4(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7) +
                                                                    to_sfixed(in_4(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8) +
                                                                    to_sfixed(in_4(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9) +
                                                                    to_sfixed(in_4(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10) +
                                                                    to_sfixed(in_4(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11) + 
                                                                    buff_1(to_integer(k_cont)), int_buff, dec_buff, fixed_saturate, fixed_truncate );
                        
                        end if;                        
                                                                    
                        temp <=    in_4(up downto down) &  
                                   in_4(up - bits downto down - bits) & 
                                   in_4(up - (bits * 2) downto down - (bits * 2)) &                         
                                   in_4(up - (bits * 3) downto down - (bits * 3)) &  
                                   in_4(up - (bits * 4) downto down - (bits * 4)) & 
                                   in_4(up - (bits * 5) downto down - (bits * 5)) & 
                                   in_4(up - (bits * 6) downto down - (bits * 6)) & 
                                   in_4(up - (bits * 7) downto down - (bits * 7)) & 
                                   in_4(up - (bits * 8) downto down - (bits * 8)) & 
                                   in_4(up - (bits * 9) downto down - (bits * 9)) & 
                                   in_4(up - (bits * 10) downto down - (bits * 10)) & 
                                   in_4(up - (bits * 11) downto down - (bits * 11));
                                   
--                             pesos(0) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)));
--                             pesos(1) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1));
--                             pesos(2) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2));
--                             pesos(3) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3));
--                             pesos(4) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4));
--                             pesos(5) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5));
--                             pesos(6) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6));
--                             pesos(7) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7));
--                             pesos(8) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8));
--                             pesos(9) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9));
--                             pesos(10) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10));
--                             pesos(11) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11));

--                             mults(0) <= resize ( to_sfixed(in_1(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(1) <= resize ( to_sfixed(in_1(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(2) <= resize ( to_sfixed(in_1(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(3) <= resize ( to_sfixed(in_1(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(4) <= resize ( to_sfixed(in_1(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(5) <= resize ( to_sfixed(in_1(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(6) <= resize ( to_sfixed(in_1(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(7) <= resize ( to_sfixed(in_1(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(8) <= resize ( to_sfixed(in_1(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(9) <= resize ( to_sfixed(in_1(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(10) <= resize ( to_sfixed(in_1(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
--                             mults(11) <= resize ( to_sfixed(in_1(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_round );
                                    
                                    
                    elsif ( (k_cont < 25) and (k_cont > 0) ) then
                    
                        k_cont <= k_cont + 1;
                        start_out <= '0';
                        pop_out <= '0';
                        
--                        pesos(0) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)));
--                             pesos(1) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1));
--                             pesos(2) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2));
--                             pesos(3) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3));
--                             pesos(4) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4));
--                             pesos(5) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5));
--                             pesos(6) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6));
--                             pesos(7) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7));
--                             pesos(8) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8));
--                             pesos(9) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9));
--                             pesos(10) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10));
--                             pesos(11) <= STD_LOGIC_VECTOR(weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11));
                             
--                         mults(0) <= resize ( to_sfixed(temp(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(1) <= resize ( to_sfixed(temp(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(2) <= resize ( to_sfixed(temp(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(3) <= resize ( to_sfixed(temp(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(4) <= resize ( to_sfixed(temp(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(5) <= resize ( to_sfixed(temp(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(6) <= resize ( to_sfixed(temp(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(7) <= resize ( to_sfixed(temp(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(8) <= resize ( to_sfixed(temp(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(9) <= resize ( to_sfixed(temp(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(10) <= resize ( to_sfixed(temp(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
--                             mults(11) <= resize ( to_sfixed(temp(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)), int_2, dec_2, fixed_saturate, fixed_truncate );
                    
                        if ( aux = 4 ) then
                        
                            buff_1(to_integer(k_cont)) <= resize (  to_sfixed(temp(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)) +
                                                                    to_sfixed(temp(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1) +
                                                                    to_sfixed(temp(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2) +
                                                                    to_sfixed(temp(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3) + 
                                                                    to_sfixed(temp(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4) +
                                                                    to_sfixed(temp(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5) +
                                                                    to_sfixed(temp(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6) +
                                                                    to_sfixed(temp(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7) +
                                                                    to_sfixed(temp(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8) +
                                                                    to_sfixed(temp(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9) +
                                                                    to_sfixed(temp(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10) +
                                                                    to_sfixed(temp(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11) + 
                                                                    buff_1(to_integer(k_cont)) + bias(to_integer(k_cont)), int_buff, dec_buff, fixed_saturate, fixed_truncate );
                                                                    
                        else
                        
                            buff_1(to_integer(k_cont)) <= resize (  to_sfixed(temp(up downto down), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12)) +
                                                                    to_sfixed(temp(up - bits downto down - bits), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 1) +
                                                                    to_sfixed(temp(up - (bits * 2) downto down - (bits * 2)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 2) +
                                                                    to_sfixed(temp(up - (bits * 3) downto down - (bits * 3)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 3) + 
                                                                    to_sfixed(temp(up - (bits * 4) downto down - (bits * 4)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 4) +
                                                                    to_sfixed(temp(up - (bits * 5) downto down - (bits * 5)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 5) +
                                                                    to_sfixed(temp(up - (bits * 6) downto down - (bits * 6)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 6) +
                                                                    to_sfixed(temp(up - (bits * 7) downto down - (bits * 7)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 7) +
                                                                    to_sfixed(temp(up - (bits * 8) downto down - (bits * 8)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 8) +
                                                                    to_sfixed(temp(up - (bits * 9) downto down - (bits * 9)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 9) +
                                                                    to_sfixed(temp(up - (bits * 10) downto down - (bits * 10)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 10) +
                                                                    to_sfixed(temp(up - (bits * 11) downto down - (bits * 11)), int_2, dec_2) * weights((to_integer(k_cont) * 60) + (to_integer(aux) * 12) + 11) + 
                                                                    buff_1(to_integer(k_cont)), int_buff, dec_buff, fixed_saturate, fixed_round );
                        
                        end if;
                                                                                                  
                    elsif (k_cont = 25 ) then
                       
                        k_cont <= "00000";
                        
                        if ( aux = 4 ) then
                        
                            aux <= "000";
                            cont <= cont + 1;
                            start_out <= '1';
                            buff_1 <= (others => X"0000");
                            
                            for i in 0 to 24 loop
                            
--                                report "capa4 " & to_hstring(STD_LOGIC_VECTOR ( buff_1(i) ));
                    
                                if ( buff_1(i) > 0 ) then
                                
                                    conv4_out((399 - (i * bits)) downto (384 - (i * bits))) <= STD_LOGIC_VECTOR ( buff_1(i) );
                                    
                                else
                                    
                                    conv4_out((399 - (i * bits)) downto (384 - (i * bits))) <= zero_out;
                                    
                                end if;
                            
                            end loop;
                        
                        else
                       
                            aux <= aux + 1;
                            start_out <= '0';
                        
                        end if;
                        
                    end if;
                    
                else
                    
                    start_out <= '0';
                    last_out <= '1';
                    
                end if;
                
            end if;

        end if;
        
    end process;
    
end Behavioral;